module Multiplier_Unit 
(
    input [6 : 0] opcode,
    input [6 : 0] funct7,
    input funct7_valid,

    input [31 : 0] bus_rs1,
    input [31 : 0] bus_rs2,

    output reg [31 : 0] mul_output
);
    
    /*

     Write your codes here
    
    */

endmodule